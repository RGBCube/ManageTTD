module main

fn main() {
	println()
}
